`ifndef WISHBONE_AGENT_TYPES_SV
  `define WISHBONE_AGENT_TYPES_SV


    typedef enum bit {WB_READ = 0, WB_WRITE = 1} wishbone_dir ;



`endif	