
`ifndef POS_L3_AGENT_PKG
  `define POS_L3_AGENT_PKG

	`include "uvm_macros.svh"
    `include "pos_l3_intf.sv"

  package pos_l3_agent_pkg;
	 import uvm_pkg::*;
	  
	  `include "pos_l3_reset_handler.sv"
	  `include "pos_l3_data_types.sv"
	  `include "pos_l3_packet.sv"
	  `include "pos_l3_agent_config.sv"
	  `include "pos_l3_item_base.sv"
      `include "pos_l3_item_drv.sv"
	  `include "pos_l3_item_mon.sv"
	  `include "pos_l3_driver.sv"
	  `include "pos_l3_sequencer.sv"
	  `include "pos_l3_monitor.sv"
	  //`include "pos_l3_coverage.sv"
	  `include "pos_l3_sequence_base.sv"
	  `include "pos_l3_sequence_simple.sv"
	  `include "pos_l3_sequence_random.sv"
	  `include "pos_l3_sequence_underflow_tx.sv"
	  `include "pos_l3_agent.sv"
	  

	 endpackage

`endif