
`ifndef POS_L3_AGENT_TYPES_SV
  `define POS_L3_AGENT_TYPES_SV

	`define LANE0        7:0
	`define LANE1       15:8
	`define LANE2      23:16
	`define LANE3      31:24
	`define LANE4      39:32
	`define LANE5      47:40
	`define LANE6      55:48
	`define LANE7      63:56
	
	`define SOP 64'h1000010000010000
	
	`define EOP 64'h00000000002c2b2a

`endif	